 `timescale 10ns / 100ps
module lesq(input [31:0]in,output [15:0]final_sqrt);
wire [31:0] data1;
wire [15:0] data2,data3,data4,data5,data6,data7;
wire odd;
wire [7:0]k,p,m;
lod ld(.in(in),.out(data1));								//find nearest power of 2^k
pe pe1(.in(data1),.out(k));									// extract value of k from 2^k
subtractor sub(.in1(in),.in2(data1),.out(data2));			//x=in-2^(k)
shifter_2 shft(.in(k),.odd(odd),.out(p));					//k/2 if k is even and (k-1)/2 if k is odd
shifter shft2(.in(data2),.in2(p),.out(data3));				//x/2^(k/2+1)
decoder de1(.in(p),.data_out(data4));						//2^(k/2)
adder add1(.in1(data3),.in2(data4),.out(data5));			//Q=2^(k/2)+x/2^(k/2+1)
error_comp ec(.in(k),.out(m));								//m-3
decoder de2(.in(m),.data_out(data6));						//2^(m-3)
adder add2(.in1(data5),.in2(data6),.out(data7));			//Q`=2^(m-3)+Q
mux mx(.in1(data7),.in2(data5),.sel(odd),.out(final_sqrt)); //ec is selected only if k is odd
endmodule


module lod(
input [31:0]in ,output reg [31:0] out
    );
    always @ (*)
	begin
	if(in[31])
	out=32'b10000000000000000000000000000000;
	else if(in[30])
	out=32'b01000000000000000000000000000000;
	else if(in[29])
	out=32'b00100000000000000000000000000000;
	else if(in[28])
	out=32'b00010000000000000000000000000000;
	else if(in[27])
	out=32'b00001000000000000000000000000000;
	else if(in[26])
	out=32'b00000100000000000000000000000000;
	else if(in[25])
	out=32'b00000010000000000000000000000000;
	else if(in[24])
	out=32'b00000001000000000000000000000000;
	else if(in[23])
	out=32'b00000000100000000000000000000000;
	else if(in[22])
	out=32'b00000000010000000000000000000000;
	else if(in[21])
	out=32'b00000000001000000000000000000000;
	else if(in[20])
	out=32'b00000000000100000000000000000000;
	else if(in[19])
	out=32'b00000000000010000000000000000000;
	else if(in[18])
	out=32'b00000000000001000000000000000000;
	else if(in[17])
	out=32'b00000000000000100000000000000000;
	else if(in[16])
	out=32'b00000000000000010000000000000000;
	else if(in[15])
	out=32'b00000000000000001000000000000000;
	else if(in[14])
	out=32'b00000000000000000100000000000000;
	else if(in[13])
	out=32'b00000000000000000010000000000000;
	else if(in[12])
	out=32'b00000000000000000001000000000000;
	else if(in[11])
	out=32'b00000000000000000000100000000000;
	else if(in[10])
	out=32'b00000000000000000000010000000000;
	else if(in[9])
	out=32'b00000000000000000000001000000000;	
	else if(in[8])
	out=32'b0000000100000000;	
    else if (in[7])
    out=32'b00000000000000000000000010000000;
    else if(in[6])
    out=32'b00000000000000000000000001000000;
    else if(in[5])
    out=32'b00000000000000000000000000100000;
    else if(in[4])
    out=32'b00000000000000000000000000010000;
    else if(in[3])
    out=32'b00000000000000000000000000001000;
    else if(in[2])
    out=32'b00000000000000000000000000000100;
    else if(in[1])
    out=32'b00000000000000000000000000000010;
	else if(in[0])
	out=32'b00000000000000000000000000000001;
    else
    out=32'b00000000000000000000000000000000;
    end
endmodule

module pe(input [31:0]in,output reg [7:0]out);
always @(*)
begin
case(in)
32'b00000000000000000000000000000001: out=8'b00000000;
32'b00000000000000000000000000000010: out=8'b00000001;
32'b00000000000000000000000000000100: out=8'b00000010;
32'b00000000000000000000000000001000: out=8'b00000011;
32'b00000000000000000000000000010000: out=8'b00000100;
32'b00000000000000000000000000100000: out=8'b00000101;
32'b00000000000000000000000001000000: out=8'b00000110;
32'b00000000000000000000000010000000: out=8'b00000111;
32'b00000000000000000000000100000000: out=8'b00001000;
32'b00000000000000000000001000000000: out=8'b00001001;
32'b00000000000000000000010000000000: out=8'b00001010;
32'b00000000000000000000100000000000: out=8'b00001011;
32'b00000000000000000001000000000000: out=8'b00001100;
32'b00000000000000000010000000000000: out=8'b00001101;
32'b00000000000000000100000000000000: out=8'b00001110;
32'b00000000000000001000000000000000: out=8'b00001111;
32'b00000000000000010000000000000000: out=8'b00010000;
32'b00000000000000100000000000000000: out=8'b00010001;
32'b00000000000001000000000000000000: out=8'b00010010;
32'b00000000000010000000000000000000: out=8'b00010011;
32'b00000000000100000000000000000000: out=8'b00010100;
32'b00000000001000000000000000000000: out=8'b00010101;
32'b00000000010000000000000000000000: out=8'b00010110;
32'b00000000100000000000000000000000: out=8'b00010111;
32'b00000001000000000000000000000000: out=8'b00011000;
32'b00000010000000000000000000000000: out=8'b00011001;
32'b00000100000000000000000000000000: out=8'b00011010;
32'b00001000000000000000000000000000: out=8'b00011011;
32'b00010000000000000000000000000000: out=8'b00011100;
32'b00100000000000000000000000000000: out=8'b00011101;
32'b01000000000000000000000000000000: out=8'b00011110;
32'b10000000000000000000000000000000: out=8'b00011111;
default: out=8'bxxxxxxxx;
endcase
end
endmodule

module subtractor(input [31:0]in1,input [31:0]in2,output [15:0]out);
reg [31:0]out1;
assign out=out1[15:0];
always@(*)
 out1=in1-in2;
endmodule



module shifter(input [15:0]in,input [7:0]in2,output [15:0]out);
reg [7:0] temp;
assign out=in>>temp;
always @(*)
temp=in2+8'b00000001;
endmodule

module shifter_2(input [7:0]in,output reg odd,output reg [7:0]out);
always @(*)
if(in[0])
begin
out=({in[7:1],1'b0})>>2'b01;
odd=1'b1;
end
else
begin
out=in>>2'b01;
odd=1'b0;
end
endmodule

module decoder(input [7:0]in,output reg [15:0]data_out);
always @(*)
case(in)
	8'b01111: data_out=16'b1000000000000000;
	8'b01110: data_out=16'b0100000000000000;
	8'b01101: data_out=16'b0010000000000000;
	8'b01100: data_out=16'b0001000000000000;
	8'b01011: data_out=16'b0000100000000000;
	8'b01010: data_out=16'b0000010000000000;
	8'b01001: data_out=16'b0000001000000000;	
	8'b01000: data_out=16'b0000000100000000;
	8'b00111: data_out=16'b0000000010000000;
	8'b00110: data_out=16'b0000000001000000;
	8'b00101: data_out=16'b0000000000100000;
	8'b00100: data_out=16'b0000000000010000;
	8'b00011: data_out=16'b0000000000001000;
	8'b00010: data_out=16'b0000000000000100;
	8'b00001: data_out=16'b0000000000000010;
	8'b00000: data_out=16'b0000000000000001;
	default: data_out=16'b0000000000000000;
endcase
endmodule

module error_comp(input [7:0]in,output reg [7:0]out);
reg [7:0]temp;
always @(*)
begin
temp=(in+8'b00000001)>>1'b1;
if(temp>=8'b00000011)
out=temp-8'b00000011;
else
out=8'b00000000;
end
endmodule

module adder(input [15:0]in1,in2,output reg [15:0]out);
always@(*)
 out=in1+in2;
endmodule

module mux(input [15:0]in1,in2,input sel,output [15:0]out);
assign out=(sel)?in1:in2;
endmodule
